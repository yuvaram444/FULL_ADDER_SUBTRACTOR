library verilog;
use verilog.vl_types.all;
entity FULL_addsub_vlg_vec_tst is
end FULL_addsub_vlg_vec_tst;
